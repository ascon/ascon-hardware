../../../LWC_rtl/FIFO.vhd