../v1/LWC_config_ccw_32.vhd