../../../LWC_rtl/PostProcessor.vhd