../v1/LWC_config_32.vhd