../../../LWC_rtl/key_piso.vhd