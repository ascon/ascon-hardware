../../../LWC_rtl/data_sipo.vhd