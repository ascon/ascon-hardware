../v1/LWC_config_ascon.vhd