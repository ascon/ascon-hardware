../v1/LWC_TB.vhd