../../../LWC_rtl/NIST_LWAPI_pkg.vhd