../../../LWC_rtl/fwft_fifo.vhd