../v1/design_pkg.vhd