../v1/CryptoCore.vhd