../../../LWC_rtl/PreProcessor.vhd